module v_telegram_bot

import net.url
