module telegram

import net.url
