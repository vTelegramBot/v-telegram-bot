/**
* Author: snxx
* For license and copyright information please follow this like:
* https://github.com/vTelegramBot/v-telegram-bot/blob/master/LICENSE
*/

module v_telegram_bot

import json


fn (bot *) send_message(c chat_table) (message, error) {
	resp, err := bot.request(c)
}

fn Bot(token string) (*bot_api, error) {
	return (token, endpoint, &http.Client{})
}

fn 
