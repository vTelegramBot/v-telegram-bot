module main
import setuper { setup }

setup(
	name='v-telegram-bot',
	version='1.0.0',
	repo='https://github.com/vTelegramBot/v-telegram-bot',
	license='MIT',
	author='snxx',
	email='snxx.lppxx@gmail.com',
	description='V for Vendetta'
)
